// jtag_to_onchipmem_32.v

// Generated using ACDS version 19.1 670

`timescale 1 ps / 1 ps
module jtag_to_onchipmem_32 (
		input  wire [13:0] avmm_pix_ram_address,    //   avmm_pix_ram.address
		input  wire        avmm_pix_ram_chipselect, //               .chipselect
		input  wire        avmm_pix_ram_clken,      //               .clken
		input  wire        avmm_pix_ram_write,      //               .write
		output wire [31:0] avmm_pix_ram_readdata,   //               .readdata
		input  wire [31:0] avmm_pix_ram_writedata,  //               .writedata
		input  wire [3:0]  avmm_pix_ram_byteenable, //               .byteenable
		input  wire        clk_clk,                 //            clk.clk
		output wire [31:0] dim_export,              //            dim.export
		output wire [31:0] hist_bins_export,        //      hist_bins.export
		input  wire [5:0]  hist_ram_address,        //       hist_ram.address
		input  wire        hist_ram_chipselect,     //               .chipselect
		input  wire        hist_ram_clken,          //               .clken
		input  wire        hist_ram_write,          //               .write
		output wire [31:0] hist_ram_readdata,       //               .readdata
		input  wire [31:0] hist_ram_writedata,      //               .writedata
		input  wire [3:0]  hist_ram_byteenable,     //               .byteenable
		output wire [31:0] mode_export,             //           mode.export
		output wire [31:0] ram_ready_export,        //      ram_ready.export
		input  wire        reset_reset_n,           //          reset.reset_n
		input  wire [31:0] start_transfer_export    // start_transfer.export
	);

	wire  [31:0] jtag_master_master_readdata;                  // mm_interconnect_0:jtag_master_master_readdata -> jtag_master:master_readdata
	wire         jtag_master_master_waitrequest;               // mm_interconnect_0:jtag_master_master_waitrequest -> jtag_master:master_waitrequest
	wire  [31:0] jtag_master_master_address;                   // jtag_master:master_address -> mm_interconnect_0:jtag_master_master_address
	wire         jtag_master_master_read;                      // jtag_master:master_read -> mm_interconnect_0:jtag_master_master_read
	wire   [3:0] jtag_master_master_byteenable;                // jtag_master:master_byteenable -> mm_interconnect_0:jtag_master_master_byteenable
	wire         jtag_master_master_readdatavalid;             // mm_interconnect_0:jtag_master_master_readdatavalid -> jtag_master:master_readdatavalid
	wire         jtag_master_master_write;                     // jtag_master:master_write -> mm_interconnect_0:jtag_master_master_write
	wire  [31:0] jtag_master_master_writedata;                 // jtag_master:master_writedata -> mm_interconnect_0:jtag_master_master_writedata
	wire         mm_interconnect_0_ram_ready_s1_chipselect;    // mm_interconnect_0:ram_ready_s1_chipselect -> ram_ready:chipselect
	wire  [31:0] mm_interconnect_0_ram_ready_s1_readdata;      // ram_ready:readdata -> mm_interconnect_0:ram_ready_s1_readdata
	wire   [1:0] mm_interconnect_0_ram_ready_s1_address;       // mm_interconnect_0:ram_ready_s1_address -> ram_ready:address
	wire         mm_interconnect_0_ram_ready_s1_write;         // mm_interconnect_0:ram_ready_s1_write -> ram_ready:write_n
	wire  [31:0] mm_interconnect_0_ram_ready_s1_writedata;     // mm_interconnect_0:ram_ready_s1_writedata -> ram_ready:writedata
	wire  [31:0] mm_interconnect_0_start_transfer_s1_readdata; // start_transfer:readdata -> mm_interconnect_0:start_transfer_s1_readdata
	wire   [1:0] mm_interconnect_0_start_transfer_s1_address;  // mm_interconnect_0:start_transfer_s1_address -> start_transfer:address
	wire         mm_interconnect_0_img_dim_s1_chipselect;      // mm_interconnect_0:img_dim_s1_chipselect -> img_dim:chipselect
	wire  [31:0] mm_interconnect_0_img_dim_s1_readdata;        // img_dim:readdata -> mm_interconnect_0:img_dim_s1_readdata
	wire   [1:0] mm_interconnect_0_img_dim_s1_address;         // mm_interconnect_0:img_dim_s1_address -> img_dim:address
	wire         mm_interconnect_0_img_dim_s1_write;           // mm_interconnect_0:img_dim_s1_write -> img_dim:write_n
	wire  [31:0] mm_interconnect_0_img_dim_s1_writedata;       // mm_interconnect_0:img_dim_s1_writedata -> img_dim:writedata
	wire         mm_interconnect_0_pixel_ram_s1_chipselect;    // mm_interconnect_0:pixel_ram_s1_chipselect -> pixel_ram:chipselect
	wire  [31:0] mm_interconnect_0_pixel_ram_s1_readdata;      // pixel_ram:readdata -> mm_interconnect_0:pixel_ram_s1_readdata
	wire  [13:0] mm_interconnect_0_pixel_ram_s1_address;       // mm_interconnect_0:pixel_ram_s1_address -> pixel_ram:address
	wire   [3:0] mm_interconnect_0_pixel_ram_s1_byteenable;    // mm_interconnect_0:pixel_ram_s1_byteenable -> pixel_ram:byteenable
	wire         mm_interconnect_0_pixel_ram_s1_write;         // mm_interconnect_0:pixel_ram_s1_write -> pixel_ram:write
	wire  [31:0] mm_interconnect_0_pixel_ram_s1_writedata;     // mm_interconnect_0:pixel_ram_s1_writedata -> pixel_ram:writedata
	wire         mm_interconnect_0_pixel_ram_s1_clken;         // mm_interconnect_0:pixel_ram_s1_clken -> pixel_ram:clken
	wire         mm_interconnect_0_hist_ram_s1_chipselect;     // mm_interconnect_0:hist_ram_s1_chipselect -> hist_ram:chipselect
	wire  [31:0] mm_interconnect_0_hist_ram_s1_readdata;       // hist_ram:readdata -> mm_interconnect_0:hist_ram_s1_readdata
	wire   [5:0] mm_interconnect_0_hist_ram_s1_address;        // mm_interconnect_0:hist_ram_s1_address -> hist_ram:address
	wire   [3:0] mm_interconnect_0_hist_ram_s1_byteenable;     // mm_interconnect_0:hist_ram_s1_byteenable -> hist_ram:byteenable
	wire         mm_interconnect_0_hist_ram_s1_write;          // mm_interconnect_0:hist_ram_s1_write -> hist_ram:write
	wire  [31:0] mm_interconnect_0_hist_ram_s1_writedata;      // mm_interconnect_0:hist_ram_s1_writedata -> hist_ram:writedata
	wire         mm_interconnect_0_hist_ram_s1_clken;          // mm_interconnect_0:hist_ram_s1_clken -> hist_ram:clken
	wire         mm_interconnect_0_mode_s1_chipselect;         // mm_interconnect_0:mode_s1_chipselect -> mode:chipselect
	wire  [31:0] mm_interconnect_0_mode_s1_readdata;           // mode:readdata -> mm_interconnect_0:mode_s1_readdata
	wire   [1:0] mm_interconnect_0_mode_s1_address;            // mm_interconnect_0:mode_s1_address -> mode:address
	wire         mm_interconnect_0_mode_s1_write;              // mm_interconnect_0:mode_s1_write -> mode:write_n
	wire  [31:0] mm_interconnect_0_mode_s1_writedata;          // mm_interconnect_0:mode_s1_writedata -> mode:writedata
	wire         mm_interconnect_0_hist_bins_s1_chipselect;    // mm_interconnect_0:hist_bins_s1_chipselect -> hist_bins:chipselect
	wire  [31:0] mm_interconnect_0_hist_bins_s1_readdata;      // hist_bins:readdata -> mm_interconnect_0:hist_bins_s1_readdata
	wire   [1:0] mm_interconnect_0_hist_bins_s1_address;       // mm_interconnect_0:hist_bins_s1_address -> hist_bins:address
	wire         mm_interconnect_0_hist_bins_s1_write;         // mm_interconnect_0:hist_bins_s1_write -> hist_bins:write_n
	wire  [31:0] mm_interconnect_0_hist_bins_s1_writedata;     // mm_interconnect_0:hist_bins_s1_writedata -> hist_bins:writedata
	wire         rst_controller_reset_out_reset;               // rst_controller:reset_out -> [hist_bins:reset_n, hist_ram:reset, hist_ram:reset2, img_dim:reset_n, mm_interconnect_0:ram_ready_reset_reset_bridge_in_reset_reset, mode:reset_n, pixel_ram:reset, pixel_ram:reset2, ram_ready:reset_n, rst_translator:in_reset, start_transfer:reset_n]
	wire         rst_controller_reset_out_reset_req;           // rst_controller:reset_req -> [hist_ram:reset_req, hist_ram:reset_req2, pixel_ram:reset_req, pixel_ram:reset_req2, rst_translator:reset_req_in]
	wire         jtag_master_master_reset_reset;               // jtag_master:master_reset_reset -> rst_controller:reset_in1
	wire         rst_controller_001_reset_out_reset;           // rst_controller_001:reset_out -> [mm_interconnect_0:jtag_master_clk_reset_reset_bridge_in_reset_reset, mm_interconnect_0:jtag_master_master_translator_reset_reset_bridge_in_reset_reset]

	jtag_to_onchipmem_32_hist_bins hist_bins (
		.clk        (clk_clk),                                   //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),           //               reset.reset_n
		.address    (mm_interconnect_0_hist_bins_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_hist_bins_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_hist_bins_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_hist_bins_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_hist_bins_s1_readdata),   //                    .readdata
		.out_port   (hist_bins_export)                           // external_connection.export
	);

	jtag_to_onchipmem_32_hist_ram hist_ram (
		.clk         (clk_clk),                                  //   clk1.clk
		.address     (mm_interconnect_0_hist_ram_s1_address),    //     s1.address
		.clken       (mm_interconnect_0_hist_ram_s1_clken),      //       .clken
		.chipselect  (mm_interconnect_0_hist_ram_s1_chipselect), //       .chipselect
		.write       (mm_interconnect_0_hist_ram_s1_write),      //       .write
		.readdata    (mm_interconnect_0_hist_ram_s1_readdata),   //       .readdata
		.writedata   (mm_interconnect_0_hist_ram_s1_writedata),  //       .writedata
		.byteenable  (mm_interconnect_0_hist_ram_s1_byteenable), //       .byteenable
		.reset       (rst_controller_reset_out_reset),           // reset1.reset
		.reset_req   (rst_controller_reset_out_reset_req),       //       .reset_req
		.address2    (hist_ram_address),                         //     s2.address
		.chipselect2 (hist_ram_chipselect),                      //       .chipselect
		.clken2      (hist_ram_clken),                           //       .clken
		.write2      (hist_ram_write),                           //       .write
		.readdata2   (hist_ram_readdata),                        //       .readdata
		.writedata2  (hist_ram_writedata),                       //       .writedata
		.byteenable2 (hist_ram_byteenable),                      //       .byteenable
		.clk2        (clk_clk),                                  //   clk2.clk
		.reset2      (rst_controller_reset_out_reset),           // reset2.reset
		.reset_req2  (rst_controller_reset_out_reset_req),       //       .reset_req
		.freeze      (1'b0)                                      // (terminated)
	);

	jtag_to_onchipmem_32_hist_bins img_dim (
		.clk        (clk_clk),                                 //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),         //               reset.reset_n
		.address    (mm_interconnect_0_img_dim_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_img_dim_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_img_dim_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_img_dim_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_img_dim_s1_readdata),   //                    .readdata
		.out_port   (dim_export)                               // external_connection.export
	);

	jtag_to_onchipmem_32_jtag_master #(
		.USE_PLI     (0),
		.PLI_PORT    (50000),
		.FIFO_DEPTHS (2)
	) jtag_master (
		.clk_clk              (clk_clk),                          //          clk.clk
		.clk_reset_reset      (~reset_reset_n),                   //    clk_reset.reset
		.master_address       (jtag_master_master_address),       //       master.address
		.master_readdata      (jtag_master_master_readdata),      //             .readdata
		.master_read          (jtag_master_master_read),          //             .read
		.master_write         (jtag_master_master_write),         //             .write
		.master_writedata     (jtag_master_master_writedata),     //             .writedata
		.master_waitrequest   (jtag_master_master_waitrequest),   //             .waitrequest
		.master_readdatavalid (jtag_master_master_readdatavalid), //             .readdatavalid
		.master_byteenable    (jtag_master_master_byteenable),    //             .byteenable
		.master_reset_reset   (jtag_master_master_reset_reset)    // master_reset.reset
	);

	jtag_to_onchipmem_32_hist_bins mode (
		.clk        (clk_clk),                              //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),      //               reset.reset_n
		.address    (mm_interconnect_0_mode_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_mode_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_mode_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_mode_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_mode_s1_readdata),   //                    .readdata
		.out_port   (mode_export)                           // external_connection.export
	);

	jtag_to_onchipmem_32_pixel_ram pixel_ram (
		.clk         (clk_clk),                                   //   clk1.clk
		.address     (mm_interconnect_0_pixel_ram_s1_address),    //     s1.address
		.clken       (mm_interconnect_0_pixel_ram_s1_clken),      //       .clken
		.chipselect  (mm_interconnect_0_pixel_ram_s1_chipselect), //       .chipselect
		.write       (mm_interconnect_0_pixel_ram_s1_write),      //       .write
		.readdata    (mm_interconnect_0_pixel_ram_s1_readdata),   //       .readdata
		.writedata   (mm_interconnect_0_pixel_ram_s1_writedata),  //       .writedata
		.byteenable  (mm_interconnect_0_pixel_ram_s1_byteenable), //       .byteenable
		.reset       (rst_controller_reset_out_reset),            // reset1.reset
		.reset_req   (rst_controller_reset_out_reset_req),        //       .reset_req
		.address2    (avmm_pix_ram_address),                      //     s2.address
		.chipselect2 (avmm_pix_ram_chipselect),                   //       .chipselect
		.clken2      (avmm_pix_ram_clken),                        //       .clken
		.write2      (avmm_pix_ram_write),                        //       .write
		.readdata2   (avmm_pix_ram_readdata),                     //       .readdata
		.writedata2  (avmm_pix_ram_writedata),                    //       .writedata
		.byteenable2 (avmm_pix_ram_byteenable),                   //       .byteenable
		.clk2        (clk_clk),                                   //   clk2.clk
		.reset2      (rst_controller_reset_out_reset),            // reset2.reset
		.reset_req2  (rst_controller_reset_out_reset_req),        //       .reset_req
		.freeze      (1'b0)                                       // (terminated)
	);

	jtag_to_onchipmem_32_hist_bins ram_ready (
		.clk        (clk_clk),                                   //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),           //               reset.reset_n
		.address    (mm_interconnect_0_ram_ready_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_ram_ready_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_ram_ready_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_ram_ready_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_ram_ready_s1_readdata),   //                    .readdata
		.out_port   (ram_ready_export)                           // external_connection.export
	);

	jtag_to_onchipmem_32_start_transfer start_transfer (
		.clk      (clk_clk),                                      //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),              //               reset.reset_n
		.address  (mm_interconnect_0_start_transfer_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_start_transfer_s1_readdata), //                    .readdata
		.in_port  (start_transfer_export)                         // external_connection.export
	);

	jtag_to_onchipmem_32_mm_interconnect_0 mm_interconnect_0 (
		.clk_src_clk_clk                                                 (clk_clk),                                      //                                               clk_src_clk.clk
		.jtag_master_clk_reset_reset_bridge_in_reset_reset               (rst_controller_001_reset_out_reset),           //               jtag_master_clk_reset_reset_bridge_in_reset.reset
		.jtag_master_master_translator_reset_reset_bridge_in_reset_reset (rst_controller_001_reset_out_reset),           // jtag_master_master_translator_reset_reset_bridge_in_reset.reset
		.ram_ready_reset_reset_bridge_in_reset_reset                     (rst_controller_reset_out_reset),               //                     ram_ready_reset_reset_bridge_in_reset.reset
		.jtag_master_master_address                                      (jtag_master_master_address),                   //                                        jtag_master_master.address
		.jtag_master_master_waitrequest                                  (jtag_master_master_waitrequest),               //                                                          .waitrequest
		.jtag_master_master_byteenable                                   (jtag_master_master_byteenable),                //                                                          .byteenable
		.jtag_master_master_read                                         (jtag_master_master_read),                      //                                                          .read
		.jtag_master_master_readdata                                     (jtag_master_master_readdata),                  //                                                          .readdata
		.jtag_master_master_readdatavalid                                (jtag_master_master_readdatavalid),             //                                                          .readdatavalid
		.jtag_master_master_write                                        (jtag_master_master_write),                     //                                                          .write
		.jtag_master_master_writedata                                    (jtag_master_master_writedata),                 //                                                          .writedata
		.hist_bins_s1_address                                            (mm_interconnect_0_hist_bins_s1_address),       //                                              hist_bins_s1.address
		.hist_bins_s1_write                                              (mm_interconnect_0_hist_bins_s1_write),         //                                                          .write
		.hist_bins_s1_readdata                                           (mm_interconnect_0_hist_bins_s1_readdata),      //                                                          .readdata
		.hist_bins_s1_writedata                                          (mm_interconnect_0_hist_bins_s1_writedata),     //                                                          .writedata
		.hist_bins_s1_chipselect                                         (mm_interconnect_0_hist_bins_s1_chipselect),    //                                                          .chipselect
		.hist_ram_s1_address                                             (mm_interconnect_0_hist_ram_s1_address),        //                                               hist_ram_s1.address
		.hist_ram_s1_write                                               (mm_interconnect_0_hist_ram_s1_write),          //                                                          .write
		.hist_ram_s1_readdata                                            (mm_interconnect_0_hist_ram_s1_readdata),       //                                                          .readdata
		.hist_ram_s1_writedata                                           (mm_interconnect_0_hist_ram_s1_writedata),      //                                                          .writedata
		.hist_ram_s1_byteenable                                          (mm_interconnect_0_hist_ram_s1_byteenable),     //                                                          .byteenable
		.hist_ram_s1_chipselect                                          (mm_interconnect_0_hist_ram_s1_chipselect),     //                                                          .chipselect
		.hist_ram_s1_clken                                               (mm_interconnect_0_hist_ram_s1_clken),          //                                                          .clken
		.img_dim_s1_address                                              (mm_interconnect_0_img_dim_s1_address),         //                                                img_dim_s1.address
		.img_dim_s1_write                                                (mm_interconnect_0_img_dim_s1_write),           //                                                          .write
		.img_dim_s1_readdata                                             (mm_interconnect_0_img_dim_s1_readdata),        //                                                          .readdata
		.img_dim_s1_writedata                                            (mm_interconnect_0_img_dim_s1_writedata),       //                                                          .writedata
		.img_dim_s1_chipselect                                           (mm_interconnect_0_img_dim_s1_chipselect),      //                                                          .chipselect
		.mode_s1_address                                                 (mm_interconnect_0_mode_s1_address),            //                                                   mode_s1.address
		.mode_s1_write                                                   (mm_interconnect_0_mode_s1_write),              //                                                          .write
		.mode_s1_readdata                                                (mm_interconnect_0_mode_s1_readdata),           //                                                          .readdata
		.mode_s1_writedata                                               (mm_interconnect_0_mode_s1_writedata),          //                                                          .writedata
		.mode_s1_chipselect                                              (mm_interconnect_0_mode_s1_chipselect),         //                                                          .chipselect
		.pixel_ram_s1_address                                            (mm_interconnect_0_pixel_ram_s1_address),       //                                              pixel_ram_s1.address
		.pixel_ram_s1_write                                              (mm_interconnect_0_pixel_ram_s1_write),         //                                                          .write
		.pixel_ram_s1_readdata                                           (mm_interconnect_0_pixel_ram_s1_readdata),      //                                                          .readdata
		.pixel_ram_s1_writedata                                          (mm_interconnect_0_pixel_ram_s1_writedata),     //                                                          .writedata
		.pixel_ram_s1_byteenable                                         (mm_interconnect_0_pixel_ram_s1_byteenable),    //                                                          .byteenable
		.pixel_ram_s1_chipselect                                         (mm_interconnect_0_pixel_ram_s1_chipselect),    //                                                          .chipselect
		.pixel_ram_s1_clken                                              (mm_interconnect_0_pixel_ram_s1_clken),         //                                                          .clken
		.ram_ready_s1_address                                            (mm_interconnect_0_ram_ready_s1_address),       //                                              ram_ready_s1.address
		.ram_ready_s1_write                                              (mm_interconnect_0_ram_ready_s1_write),         //                                                          .write
		.ram_ready_s1_readdata                                           (mm_interconnect_0_ram_ready_s1_readdata),      //                                                          .readdata
		.ram_ready_s1_writedata                                          (mm_interconnect_0_ram_ready_s1_writedata),     //                                                          .writedata
		.ram_ready_s1_chipselect                                         (mm_interconnect_0_ram_ready_s1_chipselect),    //                                                          .chipselect
		.start_transfer_s1_address                                       (mm_interconnect_0_start_transfer_s1_address),  //                                         start_transfer_s1.address
		.start_transfer_s1_readdata                                      (mm_interconnect_0_start_transfer_s1_readdata)  //                                                          .readdata
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.reset_in1      (jtag_master_master_reset_reset),     // reset_in1.reset
		.clk            (clk_clk),                            //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.clk            (clk_clk),                            //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
